m9k2_inst : m9k2 PORT MAP (
		address	 => address_sig,
		clken	 => clken_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
