/*
 *  8 bit pwm DAC
 *  Copyright (C) 2010  Donna Polehn <dpolehn@verizon.net>
 *
 *  This file is part of the Zet processor. This processor is free
 *  hardware; you can redistribute it and/or modify it under the terms of
 *  the GNU General Public License as published by the Free Software
 *  Foundation; either version 3, or (at your option) any later version.
 *
 *  Zet is distrubuted in the hope that it will be useful, but WITHOUT
 *  ANY WARRANTY; without even the implied warranty of MERCHANTABILITY
 *  or FITNESS FOR A PARTICULAR PURPOSE. See the GNU General Public
 *  License for more details.
 *
 *  You should have received a copy of the GNU General Public License
 *  along with Zet; see the file COPYING. If not, see
 *  <http://www.gnu.org/licenses/>.
 */

module sound_dac8 (
    input        clk,
    input  [7:0] dac_in,
    input        speaker,
    output       audio_out
  );

  reg [9:0] dac_register;

  assign audio_out = dac_register[9];

  always @(posedge clk) dac_register <= dac_register[7:0] + dac_in + {speaker,7'b0000000};

endmodule
