--+-----------------------------------+-------------------------------------+--
--|                      ___   ___    | (c) 2013-2014 William R Sowerbutts  |--
--|   ___  ___   ___ ___( _ ) / _ \   | will@sowerbutts.com                 |--
--|  / __|/ _ \ / __|_  / _ \| | | |  |                                     |--
--|  \__ \ (_) | (__ / / (_) | |_| |  | A Z80 FPGA computer, just for fun   |--
--|  |___/\___/ \___/___\___/ \___/   |                                     |--
--|                                   |              http://sowerbutts.com/ |--
--+-----------------------------------+-------------------------------------+--
--| An inferrable 4KB ROM to contain the monitor program                    |--
--+-------------------------------------------------------------------------+--
--
-- MonZ80_template.vhd contains the template VHDL for the ROM but no actual
-- data. The "ROMHERE" string is replaced by byte data by the "make_vhdl_rom"
-- tool in software/tools which is invoked to generate "MonZ80.vhd" after
-- the monitor program has been assembled.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity MonZ80 is
   port(
      clk           : in  std_logic;
      a             : in  std_logic_vector(11 downto 0);
      d             : out std_logic_vector(7 downto 0)
   );
end MonZ80;

architecture arch of MonZ80 is
   constant byte_rom_WIDTH: integer := 8;
   type byte_rom_type is array (0 to 4095) of std_logic_vector(byte_rom_WIDTH-1 downto 0);
   signal address_latch : std_logic_vector(11 downto 0) := (others => '0');

   -- actually memory cells
   signal byte_rom : byte_rom_type := (
   -- ROM contents follows


X"DB", X"20", X"47", X"F3", X"3E", X"0F", X"D3", X"F8", X"3E", X"20", X"D3", X"FC", X"AF", X"D3", X"FD", X"3E",
X"03", X"D3", X"FB", X"3E", X"0E", X"D3", X"F8", X"3E", X"20", X"D3", X"FC", X"3E", X"01", X"D3", X"FD", X"3E",
X"03", X"D3", X"FB", X"C3", X"26", X"F0", X"AF", X"D3", X"F8", X"D3", X"FC", X"D3", X"FD", X"3E", X"03", X"D3",
X"FB", X"78", X"31", X"00", X"F0", X"21", X"27", X"F7", X"CD", X"0B", X"F6", X"21", X"00", X"00", X"3E", X"01",
X"D3", X"F8", X"3E", X"03", X"D3", X"FB", X"7C", X"D3", X"FC", X"D3", X"21", X"7D", X"D3", X"FD", X"E5", X"21",
X"00", X"10", X"11", X"01", X"10", X"01", X"FF", X"0F", X"36", X"00", X"ED", X"B0", X"E1", X"23", X"7D", X"FE",
X"00", X"20", X"E3", X"7C", X"CD", X"57", X"F6", X"7C", X"FE", X"08", X"20", X"DA", X"CD", X"22", X"F6", X"AF",
X"D3", X"21", X"AF", X"D3", X"FC", X"3C", X"D3", X"FD", X"31", X"00", X"F0", X"FD", X"21", X"00", X"EF", X"3E",
X"C3", X"32", X"00", X"00", X"21", X"26", X"F0", X"22", X"01", X"00", X"AF", X"D3", X"21", X"21", X"41", X"F7",
X"CD", X"0B", X"F6", X"DB", X"01", X"DB", X"00", X"CB", X"7F", X"20", X"F8", X"21", X"17", X"F8", X"CD", X"0B",
X"F6", X"FD", X"E5", X"E1", X"CD", X"72", X"F6", X"CD", X"22", X"F6", X"DD", X"21", X"5F", X"FD", X"FD", X"E5",
X"E1", X"7E", X"FE", X"00", X"28", X"E5", X"DD", X"5E", X"00", X"DD", X"56", X"01", X"CD", X"01", X"F6", X"CA",
X"D9", X"F0", X"01", X"04", X"00", X"DD", X"09", X"DD", X"7E", X"00", X"DD", X"B6", X"01", X"FE", X"00", X"20",
X"DD", X"21", X"1D", X"F8", X"CD", X"0B", X"F6", X"18", X"C2", X"DD", X"5E", X"02", X"DD", X"56", X"03", X"D5",
X"DD", X"E1", X"DD", X"E9", X"21", X"42", X"FA", X"CD", X"0B", X"F6", X"C3", X"9B", X"F0", X"CD", X"EF", X"F6",
X"CD", X"FF", X"F6", X"D5", X"CD", X"3F", X"F6", X"3E", X"3D", X"CD", X"65", X"F6", X"3E", X"20", X"CD", X"65",
X"F6", X"C1", X"ED", X"78", X"CD", X"48", X"F6", X"CD", X"22", X"F6", X"CD", X"EF", X"F6", X"7E", X"FE", X"00",
X"CA", X"9B", X"F0", X"18", X"D8", X"CD", X"EF", X"F6", X"CD", X"FF", X"F6", X"D5", X"CD", X"EF", X"F6", X"CD",
X"FF", X"F6", X"7A", X"FE", X"00", X"20", X"31", X"C1", X"ED", X"59", X"03", X"CD", X"EF", X"F6", X"7E", X"FE",
X"00", X"CA", X"9B", X"F0", X"C5", X"18", X"E5", X"CD", X"EF", X"F6", X"CD", X"FF", X"F6", X"D5", X"DD", X"E1",
X"CD", X"EF", X"F6", X"7E", X"FE", X"00", X"CA", X"9B", X"F0", X"CD", X"05", X"F7", X"7A", X"FE", X"00", X"20",
X"07", X"DD", X"73", X"00", X"DD", X"23", X"18", X"E8", X"21", X"5A", X"F8", X"CD", X"0B", X"F6", X"C3", X"9B",
X"F0", X"CD", X"EF", X"F6", X"CD", X"FF", X"F6", X"D5", X"CD", X"EF", X"F6", X"CD", X"05", X"F7", X"7B", X"B2",
X"FE", X"00", X"20", X"02", X"1E", X"01", X"E1", X"CD", X"7D", X"F1", X"C3", X"9B", X"F0", X"CD", X"2D", X"F6",
X"3E", X"3A", X"CD", X"65", X"F6", X"3E", X"20", X"CD", X"65", X"F6", X"7E", X"CD", X"48", X"F6", X"23", X"1B",
X"7B", X"B2", X"28", X"0C", X"7D", X"E6", X"0F", X"FE", X"00", X"20", X"EA", X"CD", X"22", X"F6", X"18", X"DD",
X"CD", X"22", X"F6", X"C9", X"CD", X"EF", X"F6", X"CD", X"FF", X"F6", X"EB", X"01", X"78", X"F0", X"C5", X"E9",
X"CD", X"EF", X"F6", X"CD", X"FF", X"F6", X"D5", X"3E", X"FF", X"D3", X"F8", X"7A", X"06", X"04", X"CB", X"3F",
X"10", X"FC", X"D3", X"FC", X"06", X"04", X"7A", X"4B", X"CB", X"21", X"17", X"10", X"FB", X"D3", X"FD", X"79",
X"F6", X"0F", X"D3", X"FE", X"3E", X"FC", X"D3", X"FF", X"DB", X"FA", X"FE", X"BA", X"20", X"31", X"DB", X"FA",
X"FE", X"BE", X"20", X"2B", X"DB", X"FA", X"6F", X"DB", X"FA", X"67", X"79", X"D3", X"FE", X"AF", X"D3", X"FF",
X"E5", X"21", X"F8", X"F8", X"CD", X"0B", X"F6", X"E1", X"E5", X"CD", X"2D", X"F6", X"CD", X"22", X"F6", X"0E",
X"FA", X"16", X"10", X"06", X"00", X"ED", X"B2", X"15", X"20", X"FB", X"DD", X"E1", X"E1", X"DD", X"E9", X"21",
X"24", X"F9", X"CD", X"0B", X"F6", X"C3", X"9B", X"F0", X"21", X"A6", X"F8", X"CD", X"0B", X"F6", X"DB", X"F8",
X"F5", X"1E", X"00", X"7B", X"D3", X"F8", X"07", X"07", X"07", X"07", X"57", X"CD", X"48", X"F6", X"3E", X"00",
X"CD", X"48", X"F6", X"3E", X"2D", X"CD", X"65", X"F6", X"7A", X"F6", X"0F", X"CD", X"48", X"F6", X"3E", X"FF",
X"CD", X"48", X"F6", X"3E", X"09", X"CD", X"65", X"F6", X"DB", X"FC", X"CD", X"48", X"F6", X"DB", X"FD", X"CD",
X"48", X"F6", X"3E", X"00", X"CD", X"48", X"F6", X"3E", X"30", X"CD", X"65", X"F6", X"3E", X"2D", X"CD", X"65",
X"F6", X"DB", X"FC", X"CD", X"48", X"F6", X"DB", X"FD", X"CD", X"48", X"F6", X"3E", X"FF", X"CD", X"48", X"F6",
X"3E", X"46", X"CD", X"65", X"F6", X"3E", X"09", X"CD", X"65", X"F6", X"3E", X"09", X"CD", X"65", X"F6", X"DB",
X"FB", X"57", X"CD", X"48", X"F6", X"3E", X"20", X"CD", X"65", X"F6", X"7A", X"E6", X"02", X"28", X"06", X"21",
X"D7", X"F8", X"CD", X"0B", X"F6", X"7A", X"E6", X"01", X"28", X"06", X"21", X"D1", X"F8", X"CD", X"0B", X"F6",
X"CD", X"22", X"F6", X"1C", X"7B", X"FE", X"10", X"C2", X"23", X"F2", X"21", X"DE", X"F8", X"CD", X"0B", X"F6",
X"3E", X"FF", X"D3", X"F8", X"DB", X"FC", X"CD", X"48", X"F6", X"DB", X"FD", X"CD", X"48", X"F6", X"DB", X"FE",
X"CD", X"48", X"F6", X"DB", X"FF", X"CD", X"48", X"F6", X"CD", X"22", X"F6", X"F1", X"D3", X"F8", X"C3", X"9B",
X"F0", X"CD", X"EF", X"F6", X"CD", X"FF", X"F6", X"D5", X"CD", X"EF", X"F6", X"CD", X"FF", X"F6", X"D5", X"CD",
X"EF", X"F6", X"CD", X"FF", X"F6", X"D5", X"C1", X"D1", X"E1", X"ED", X"B0", X"C3", X"9B", X"F0", X"CD", X"EF",
X"F6", X"7E", X"FE", X"00", X"28", X"06", X"CD", X"05", X"F7", X"D5", X"E1", X"F9", X"21", X"60", X"F9", X"CD",
X"0B", X"F6", X"21", X"00", X"00", X"39", X"CD", X"2D", X"F6", X"CD", X"22", X"F6", X"C3", X"9B", X"F0", X"CD",
X"EF", X"F6", X"7E", X"FE", X"00", X"28", X"06", X"CD", X"05", X"F7", X"D5", X"FD", X"E1", X"21", X"64", X"F9",
X"CD", X"0B", X"F6", X"FD", X"E5", X"E1", X"CD", X"2D", X"F6", X"CD", X"22", X"F6", X"C3", X"9B", X"F0", X"CD",
X"EF", X"F6", X"11", X"00", X"02", X"7E", X"FE", X"00", X"28", X"03", X"CD", X"05", X"F7", X"21", X"97", X"F9",
X"CD", X"0B", X"F6", X"CD", X"3F", X"F6", X"CD", X"9C", X"F3", X"3E", X"0D", X"D3", X"F8", X"DB", X"FC", X"47",
X"DB", X"FD", X"4F", X"C5", X"CD", X"22", X"F6", X"01", X"00", X"02", X"EB", X"CD", X"2D", X"F6", X"7D", X"E6",
X"0F", X"FE", X"0F", X"20", X"05", X"CD", X"22", X"F6", X"18", X"05", X"3E", X"20", X"CD", X"65", X"F6", X"7C",
X"D3", X"FC", X"7D", X"D3", X"FD", X"E5", X"C5", X"21", X"00", X"D0", X"11", X"01", X"D0", X"01", X"FF", X"0F",
X"3E", X"E5", X"77", X"ED", X"B0", X"C1", X"E1", X"23", X"0B", X"78", X"B1", X"FE", X"00", X"20", X"CC", X"CD",
X"22", X"F6", X"C1", X"78", X"D3", X"FC", X"79", X"D3", X"FD", X"C3", X"9B", X"F0", X"21", X"1B", X"FA", X"CD",
X"0B", X"F6", X"CD", X"E6", X"F6", X"E6", X"DF", X"FE", X"59", X"C8", X"FE", X"4E", X"20", X"F4", X"CD", X"22",
X"F6", X"E1", X"C3", X"9B", X"F0", X"E5", X"CD", X"74", X"F5", X"E1", X"CD", X"EF", X"F6", X"01", X"00", X"02",
X"11", X"00", X"02", X"7E", X"FE", X"00", X"28", X"1A", X"CD", X"05", X"F7", X"CD", X"EF", X"F6", X"7E", X"FE",
X"00", X"28", X"0F", X"D5", X"CD", X"05", X"F7", X"7A", X"E6", X"F0", X"FE", X"00", X"C2", X"58", X"F1", X"D5",
X"C1", X"D1", X"21", X"B8", X"F9", X"CD", X"0B", X"F6", X"CD", X"3F", X"F6", X"21", X"D8", X"F9", X"CD", X"0B",
X"F6", X"CD", X"36", X"F6", X"CD", X"9C", X"F3", X"CD", X"22", X"F6", X"3E", X"04", X"A7", X"CB", X"11", X"CB",
X"10", X"3D", X"FE", X"00", X"20", X"F6", X"3E", X"0D", X"D3", X"F8", X"DB", X"FC", X"67", X"DB", X"FD", X"6F",
X"E5", X"C5", X"E1", X"01", X"00", X"02", X"CD", X"3F", X"F6", X"7B", X"E6", X"0F", X"FE", X"0F", X"20", X"05",
X"CD", X"22", X"F6", X"18", X"05", X"3E", X"20", X"CD", X"65", X"F6", X"7A", X"D3", X"FC", X"7B", X"D3", X"FD",
X"D5", X"E5", X"CD", X"CC", X"F5", X"3E", X"0B", X"D3", X"1A", X"CD", X"61", X"F4", X"D3", X"1A", X"21", X"00",
X"D0", X"D3", X"1A", X"DB", X"1B", X"77", X"23", X"7C", X"FE", X"E0", X"20", X"F5", X"CD", X"C7", X"F5", X"E1",
X"11", X"10", X"00", X"19", X"D1", X"13", X"0B", X"78", X"B1", X"20", X"BB", X"CD", X"22", X"F6", X"C3", X"92",
X"F3", X"7C", X"D3", X"1A", X"7D", X"D3", X"1A", X"AF", X"D3", X"1A", X"C9", X"E5", X"CD", X"74", X"F5", X"E1",
X"CD", X"EF", X"F6", X"01", X"00", X"02", X"11", X"00", X"02", X"7E", X"FE", X"00", X"28", X"1A", X"CD", X"05",
X"F7", X"CD", X"EF", X"F6", X"7E", X"FE", X"00", X"28", X"0F", X"D5", X"CD", X"05", X"F7", X"7A", X"E6", X"F0",
X"FE", X"00", X"C2", X"58", X"F1", X"D5", X"C1", X"D1", X"21", X"EA", X"F9", X"CD", X"0B", X"F6", X"CD", X"3F",
X"F6", X"21", X"0B", X"FA", X"CD", X"0B", X"F6", X"CD", X"36", X"F6", X"CD", X"9C", X"F3", X"CD", X"22", X"F6",
X"3E", X"04", X"A7", X"CB", X"11", X"CB", X"10", X"3D", X"FE", X"00", X"20", X"F6", X"3E", X"0D", X"D3", X"F8",
X"DB", X"FC", X"67", X"DB", X"FD", X"6F", X"E5", X"C5", X"E1", X"01", X"00", X"02", X"CD", X"3F", X"F6", X"7B",
X"E6", X"0F", X"FE", X"0F", X"20", X"05", X"CD", X"22", X"F6", X"18", X"05", X"3E", X"20", X"CD", X"65", X"F6",
X"D5", X"7A", X"D3", X"FC", X"7B", X"D3", X"FD", X"CD", X"49", X"F5", X"FE", X"00", X"28", X"4A", X"E5", X"CD",
X"F2", X"F5", X"CD", X"CC", X"F5", X"3E", X"20", X"D3", X"1A", X"CD", X"61", X"F4", X"CD", X"C7", X"F5", X"11",
X"00", X"D0", X"CD", X"F2", X"F5", X"CD", X"CC", X"F5", X"3E", X"02", X"D3", X"1A", X"CD", X"61", X"F4", X"1A",
X"D3", X"1A", X"13", X"7B", X"FE", X"00", X"20", X"F7", X"CD", X"C7", X"F5", X"23", X"7A", X"FE", X"E0", X"20",
X"E1", X"E1", X"CD", X"EA", X"F5", X"CD", X"49", X"F5", X"FE", X"00", X"28", X"0C", X"CD", X"22", X"F6", X"21",
X"23", X"FA", X"CD", X"0B", X"F6", X"CD", X"58", X"F1", X"11", X"10", X"00", X"19", X"D1", X"13", X"0B", X"78",
X"B1", X"20", X"89", X"CD", X"22", X"F6", X"C3", X"92", X"F3", X"E5", X"CD", X"CC", X"F5", X"3E", X"0B", X"D3",
X"1A", X"CD", X"61", X"F4", X"D3", X"1A", X"21", X"00", X"D0", X"D3", X"1A", X"DB", X"1B", X"BE", X"20", X"0D",
X"23", X"7C", X"FE", X"E0", X"20", X"F3", X"CD", X"C7", X"F5", X"E1", X"3E", X"00", X"C9", X"CD", X"C7", X"F5",
X"E1", X"3E", X"FF", X"C9", X"CD", X"C3", X"F5", X"21", X"69", X"F9", X"CD", X"0B", X"F6", X"CD", X"CC", X"F5",
X"3E", X"9F", X"D3", X"1A", X"AF", X"D3", X"1A", X"D3", X"1A", X"D3", X"1A", X"D3", X"1A", X"DB", X"1B", X"67",
X"D3", X"1A", X"DB", X"1B", X"6F", X"D3", X"1A", X"DB", X"1B", X"5F", X"CD", X"C7", X"F5", X"CD", X"2D", X"F6",
X"7B", X"CD", X"48", X"F6", X"7C", X"FE", X"C2", X"20", X"11", X"7D", X"FE", X"20", X"20", X"0C", X"7B", X"FE",
X"17", X"20", X"07", X"21", X"83", X"F9", X"CD", X"0B", X"F6", X"C9", X"21", X"8B", X"F9", X"CD", X"0B", X"F6",
X"C3", X"9B", X"F0", X"3E", X"01", X"D3", X"1C", X"3E", X"FF", X"D3", X"18", X"C9", X"3E", X"FE", X"D3", X"18",
X"C9", X"CD", X"CC", X"F5", X"3E", X"06", X"D3", X"1A", X"CD", X"C7", X"F5", X"CD", X"CC", X"F5", X"3E", X"05",
X"D3", X"1A", X"D3", X"1A", X"CD", X"C7", X"F5", X"DB", X"1B", X"C9", X"CD", X"DB", X"F5", X"CB", X"47", X"C8",
X"18", X"F8", X"CD", X"DB", X"F5", X"CB", X"47", X"20", X"F9", X"CB", X"4F", X"C0", X"CD", X"D1", X"F5", X"18",
X"F1", X"1A", X"FE", X"00", X"C8", X"BE", X"C0", X"13", X"23", X"18", X"F6", X"7E", X"A7", X"C8", X"CD", X"65",
X"F6", X"23", X"18", X"F7", X"7E", X"A7", X"C8", X"CD", X"48", X"F6", X"3E", X"20", X"CD", X"65", X"F6", X"23",
X"18", X"F2", X"3E", X"0D", X"CD", X"65", X"F6", X"3E", X"0A", X"CD", X"65", X"F6", X"C9", X"7C", X"CD", X"48",
X"F6", X"7D", X"CD", X"48", X"F6", X"C9", X"78", X"CD", X"48", X"F6", X"79", X"CD", X"48", X"F6", X"C9", X"7A",
X"CD", X"48", X"F6", X"7B", X"CD", X"48", X"F6", X"C9", X"C5", X"4F", X"1F", X"1F", X"1F", X"1F", X"CD", X"57",
X"F6", X"79", X"CD", X"57", X"F6", X"C1", X"C9", X"E6", X"0F", X"FE", X"0A", X"38", X"02", X"C6", X"07", X"C6",
X"30", X"CD", X"65", X"F6", X"C9", X"C5", X"47", X"DB", X"00", X"CB", X"77", X"20", X"FA", X"78", X"D3", X"01",
X"C1", X"C9", X"0E", X"00", X"CD", X"E6", X"F6", X"FE", X"40", X"20", X"08", X"CD", X"65", X"F6", X"18", X"41",
X"CD", X"E6", X"F6", X"FE", X"0D", X"28", X"36", X"FE", X"0A", X"28", X"32", X"FE", X"08", X"28", X"16", X"FE",
X"7F", X"28", X"12", X"FE", X"20", X"DA", X"80", X"F6", X"FE", X"7F", X"D2", X"80", X"F6", X"77", X"23", X"0C",
X"CD", X"65", X"F6", X"18", X"DB", X"79", X"FE", X"00", X"28", X"D6", X"2B", X"0D", X"3E", X"08", X"CD", X"65",
X"F6", X"3E", X"20", X"CD", X"65", X"F6", X"3E", X"08", X"CD", X"65", X"F6", X"18", X"C3", X"3E", X"00", X"77",
X"C9", X"CD", X"E6", X"F6", X"FE", X"0D", X"28", X"F5", X"FE", X"0A", X"28", X"F1", X"77", X"23", X"FE", X"20",
X"28", X"05", X"CD", X"65", X"F6", X"18", X"EA", X"CD", X"E6", X"F6", X"FE", X"0D", X"28", X"DF", X"FE", X"0A",
X"28", X"DB", X"77", X"23", X"18", X"F1", X"DB", X"00", X"CB", X"7F", X"28", X"FA", X"DB", X"01", X"C9", X"7E",
X"FE", X"20", X"C0", X"23", X"18", X"F9", X"FE", X"61", X"D8", X"FE", X"7B", X"D0", X"E6", X"5F", X"C9", X"7E",
X"FE", X"00", X"CA", X"58", X"F1", X"16", X"00", X"1E", X"00", X"7E", X"FE", X"30", X"D8", X"FE", X"40", X"38",
X"02", X"D6", X"07", X"D6", X"30", X"E6", X"0F", X"C5", X"06", X"04", X"A7", X"CB", X"13", X"CB", X"12", X"10",
X"F9", X"C1", X"B3", X"5F", X"23", X"18", X"E2", X"0D", X"0A", X"43", X"6F", X"6C", X"64", X"20", X"62", X"6F",
X"6F", X"74", X"3A", X"20", X"7A", X"65", X"72", X"6F", X"69", X"6E", X"67", X"20", X"52", X"41", X"4D", X"20",
X"00", X"0D", X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20",
X"20", X"20", X"20", X"20", X"20", X"20", X"5F", X"5F", X"5F", X"20", X"20", X"20", X"5F", X"5F", X"5F", X"20",
X"20", X"0D", X"0A", X"20", X"5F", X"5F", X"5F", X"20", X"20", X"5F", X"5F", X"5F", X"20", X"20", X"20", X"5F",
X"5F", X"5F", X"20", X"5F", X"5F", X"5F", X"28", X"20", X"5F", X"20", X"29", X"20", X"2F", X"20", X"5F", X"20",
X"5C", X"20", X"0D", X"0A", X"2F", X"20", X"5F", X"5F", X"7C", X"2F", X"20", X"5F", X"20", X"5C", X"20", X"2F",
X"20", X"5F", X"5F", X"7C", X"5F", X"20", X"20", X"2F", X"20", X"5F", X"20", X"5C", X"7C", X"20", X"7C", X"20",
X"7C", X"20", X"7C", X"0D", X"0A", X"5C", X"5F", X"5F", X"20", X"5C", X"20", X"28", X"5F", X"29", X"20", X"7C",
X"20", X"28", X"5F", X"5F", X"20", X"2F", X"20", X"2F", X"20", X"28", X"5F", X"29", X"20", X"7C", X"20", X"7C",
X"5F", X"7C", X"20", X"7C", X"0D", X"0A", X"7C", X"5F", X"5F", X"5F", X"2F", X"5C", X"5F", X"5F", X"5F", X"2F",
X"20", X"5C", X"5F", X"5F", X"5F", X"2F", X"5F", X"5F", X"5F", X"5C", X"5F", X"5F", X"5F", X"2F", X"20", X"5C",
X"5F", X"5F", X"5F", X"2F", X"20", X"0D", X"0A", X"5A", X"38", X"30", X"20", X"52", X"4F", X"4D", X"20", X"4D",
X"6F", X"6E", X"69", X"74", X"6F", X"72", X"20", X"28", X"57", X"69", X"6C", X"6C", X"20", X"53", X"6F", X"77",
X"65", X"72", X"62", X"75", X"74", X"74", X"73", X"2C", X"20", X"32", X"30", X"31", X"33", X"2D", X"31", X"32",
X"2D", X"31", X"32", X"29", X"0D", X"0A", X"00", X"5A", X"38", X"30", X"3E", X"20", X"00", X"45", X"72", X"72",
X"6F", X"72", X"20", X"72", X"65", X"64", X"75", X"63", X"65", X"73", X"0D", X"0A", X"59", X"6F", X"75", X"72",
X"20", X"65", X"78", X"70", X"65", X"6E", X"73", X"69", X"76", X"65", X"20", X"63", X"6F", X"6D", X"70", X"75",
X"74", X"65", X"72", X"0D", X"0A", X"54", X"6F", X"20", X"61", X"20", X"73", X"69", X"6D", X"70", X"6C", X"65",
X"20", X"73", X"74", X"6F", X"6E", X"65", X"2E", X"0D", X"0A", X"00", X"45", X"72", X"72", X"6F", X"72", X"73",
X"20", X"68", X"61", X"76", X"65", X"20", X"6F", X"63", X"63", X"75", X"72", X"72", X"65", X"64", X"2E", X"0D",
X"0A", X"57", X"65", X"20", X"77", X"6F", X"6E", X"27", X"74", X"20", X"74", X"65", X"6C", X"6C", X"20", X"79",
X"6F", X"75", X"20", X"77", X"68", X"65", X"72", X"65", X"20", X"6F", X"72", X"20", X"77", X"68", X"79", X"2E",
X"0D", X"0A", X"4C", X"61", X"7A", X"79", X"20", X"70", X"72", X"6F", X"67", X"72", X"61", X"6D", X"6D", X"65",
X"72", X"73", X"2E", X"0D", X"0A", X"00", X"56", X"69", X"72", X"74", X"75", X"61", X"6C", X"20", X"28", X"46",
X"38", X"29", X"09", X"50", X"68", X"79", X"73", X"69", X"63", X"61", X"6C", X"20", X"28", X"46", X"43", X"20",
X"46", X"44", X"29", X"09", X"46", X"6C", X"61", X"67", X"73", X"20", X"28", X"46", X"42", X"29", X"0D", X"0A",
X"00", X"52", X"45", X"41", X"44", X"20", X"00", X"57", X"52", X"49", X"54", X"45", X"20", X"00", X"31", X"37",
X"74", X"68", X"20", X"50", X"61", X"67", X"65", X"20", X"50", X"6F", X"69", X"6E", X"74", X"65", X"72", X"20",
X"28", X"46", X"41", X"29", X"20", X"3D", X"20", X"00", X"4C", X"6F", X"61", X"64", X"69", X"6E", X"67", X"20",
X"73", X"74", X"61", X"67", X"65", X"20", X"32", X"20", X"62", X"6F", X"6F", X"74", X"73", X"74", X"72", X"61",
X"70", X"20", X"66", X"72", X"6F", X"6D", X"20", X"52", X"41", X"4D", X"20", X"64", X"69", X"73", X"6B", X"20",
X"74", X"6F", X"20", X"00", X"42", X"61", X"64", X"20", X"6D", X"61", X"67", X"69", X"63", X"20", X"6E", X"75",
X"6D", X"62", X"65", X"72", X"2E", X"20", X"47", X"65", X"6E", X"74", X"6C", X"65", X"6D", X"65", X"6E", X"2C",
X"20", X"70", X"6C", X"65", X"61", X"73", X"65", X"20", X"63", X"68", X"65", X"63", X"6B", X"20", X"79", X"6F",
X"75", X"72", X"20", X"52", X"41", X"4D", X"20", X"64", X"69", X"73", X"6B", X"73", X"2E", X"0D", X"0A", X"00",
X"53", X"50", X"3D", X"00", X"42", X"55", X"46", X"3D", X"00", X"43", X"68", X"65", X"63", X"6B", X"69", X"6E",
X"67", X"20", X"53", X"50", X"49", X"20", X"66", X"6C", X"61", X"73", X"68", X"20", X"74", X"79", X"70", X"65",
X"3A", X"20", X"00", X"20", X"28", X"4F", X"4B", X"29", X"0D", X"0A", X"00", X"20", X"46", X"41", X"49", X"4C",
X"21", X"20", X"3A", X"28", X"0D", X"0A", X"00", X"45", X"72", X"61", X"73", X"65", X"20", X"52", X"41", X"4D",
X"20", X"64", X"69", X"73", X"6B", X"20", X"73", X"74", X"61", X"72", X"74", X"69", X"6E", X"67", X"20", X"61",
X"74", X"20", X"70", X"61", X"67", X"65", X"20", X"00", X"52", X"65", X"61", X"64", X"20", X"52", X"41", X"4D",
X"20", X"64", X"69", X"73", X"6B", X"20", X"73", X"74", X"61", X"72", X"74", X"69", X"6E", X"67", X"20", X"61",
X"74", X"20", X"70", X"61", X"67", X"65", X"20", X"00", X"20", X"66", X"72", X"6F", X"6D", X"20", X"66", X"6C",
X"61", X"73", X"68", X"20", X"70", X"61", X"67", X"65", X"20", X"00", X"57", X"72", X"69", X"74", X"65", X"20",
X"52", X"41", X"4D", X"20", X"64", X"69", X"73", X"6B", X"20", X"73", X"74", X"61", X"72", X"74", X"69", X"6E",
X"67", X"20", X"61", X"74", X"20", X"70", X"61", X"67", X"65", X"20", X"00", X"20", X"74", X"6F", X"20", X"66",
X"6C", X"61", X"73", X"68", X"20", X"70", X"61", X"67", X"65", X"20", X"00", X"20", X"28", X"79", X"2F", X"6E",
X"29", X"3F", X"00", X"46", X"6C", X"61", X"73", X"68", X"20", X"77", X"72", X"69", X"74", X"65", X"20", X"76",
X"65", X"72", X"69", X"66", X"79", X"20", X"66", X"61", X"69", X"6C", X"65", X"64", X"20", X"3A", X"28", X"0D",
X"0A", X"00", X"43", X"6F", X"6D", X"6D", X"61", X"6E", X"64", X"73", X"3A", X"0D", X"0A", X"09", X"64", X"6D",
X"20", X"61", X"64", X"64", X"72", X"20", X"5B", X"6C", X"65", X"6E", X"5D", X"09", X"09", X"09", X"64", X"69",
X"73", X"70", X"6C", X"61", X"79", X"20", X"6D", X"65", X"6D", X"6F", X"72", X"79", X"20", X"63", X"6F", X"6E",
X"74", X"65", X"6E", X"74", X"73", X"20", X"66", X"72", X"6F", X"6D", X"20", X"61", X"64", X"64", X"72", X"20",
X"66", X"6F", X"72", X"20", X"6C", X"65", X"6E", X"20", X"28", X"64", X"65", X"66", X"61", X"75", X"6C", X"74",
X"20", X"31", X"29", X"20", X"62", X"79", X"74", X"65", X"73", X"0D", X"0A", X"09", X"77", X"6D", X"20", X"61",
X"64", X"64", X"72", X"20", X"76", X"61", X"6C", X"20", X"5B", X"76", X"61", X"6C", X"2E", X"2E", X"2E", X"5D",
X"09", X"09", X"77", X"72", X"69", X"74", X"65", X"20", X"62", X"79", X"74", X"65", X"73", X"20", X"74", X"6F",
X"20", X"6D", X"65", X"6D", X"6F", X"72", X"79", X"20", X"73", X"74", X"61", X"72", X"74", X"69", X"6E", X"67",
X"20", X"61", X"74", X"20", X"61", X"64", X"64", X"72", X"0D", X"0A", X"09", X"63", X"70", X"20", X"73", X"72",
X"63", X"20", X"64", X"73", X"74", X"20", X"6C", X"65", X"6E", X"09", X"09", X"09", X"63", X"6F", X"70", X"79",
X"20", X"6C", X"65", X"6E", X"20", X"62", X"79", X"74", X"65", X"73", X"20", X"66", X"72", X"6F", X"6D", X"20",
X"73", X"72", X"63", X"20", X"74", X"6F", X"20", X"64", X"73", X"74", X"0D", X"0A", X"09", X"72", X"75", X"6E",
X"20", X"61", X"64", X"64", X"72", X"09", X"09", X"09", X"72", X"75", X"6E", X"20", X"63", X"6F", X"64", X"65",
X"20", X"61", X"74", X"20", X"61", X"64", X"64", X"72", X"0D", X"0A", X"09", X"69", X"6E", X"20", X"61", X"64",
X"64", X"72", X"09", X"09", X"09", X"09", X"72", X"65", X"61", X"64", X"20", X"49", X"2F", X"4F", X"20", X"70",
X"6F", X"72", X"74", X"20", X"61", X"74", X"20", X"61", X"64", X"64", X"72", X"2C", X"20", X"64", X"69", X"73",
X"70", X"6C", X"61", X"79", X"20", X"72", X"65", X"73", X"75", X"6C", X"74", X"0D", X"0A", X"09", X"6F", X"75",
X"74", X"20", X"61", X"64", X"64", X"72", X"20", X"76", X"61", X"6C", X"20", X"5B", X"76", X"61", X"6C", X"2E",
X"2E", X"2E", X"5D", X"09", X"09", X"77", X"72", X"69", X"74", X"65", X"20", X"49", X"2F", X"4F", X"20", X"70",
X"6F", X"72", X"74", X"20", X"61", X"74", X"20", X"61", X"64", X"64", X"72", X"20", X"77", X"69", X"74", X"68",
X"20", X"76", X"61", X"6C", X"0D", X"0A", X"09", X"6D", X"6D", X"75", X"09", X"09", X"09", X"09", X"73", X"68",
X"6F", X"77", X"20", X"4D", X"4D", X"55", X"20", X"73", X"74", X"61", X"74", X"65", X"0D", X"0A", X"09", X"73",
X"70", X"20", X"5B", X"61", X"64", X"64", X"72", X"5D", X"09", X"09", X"09", X"73", X"68", X"6F", X"77", X"20",
X"73", X"74", X"61", X"63", X"6B", X"20", X"70", X"6F", X"69", X"6E", X"74", X"65", X"72", X"20", X"28", X"61",
X"6E", X"64", X"20", X"73", X"65", X"74", X"20", X"74", X"6F", X"20", X"61", X"64", X"64", X"72", X"29", X"0D",
X"0A", X"09", X"62", X"75", X"66", X"20", X"5B", X"61", X"64", X"64", X"72", X"5D", X"09", X"09", X"09", X"73",
X"68", X"6F", X"77", X"20", X"69", X"6E", X"70", X"75", X"74", X"20", X"62", X"75", X"66", X"66", X"65", X"72",
X"20", X"28", X"61", X"6E", X"64", X"20", X"73", X"65", X"74", X"20", X"74", X"6F", X"20", X"61", X"64", X"64",
X"72", X"29", X"0D", X"0A", X"09", X"72", X"62", X"6F", X"6F", X"74", X"20", X"70", X"61", X"67", X"65", X"09",
X"09", X"09", X"42", X"6F", X"6F", X"74", X"20", X"66", X"72", X"6F", X"6D", X"20", X"52", X"41", X"4D", X"20",
X"64", X"69", X"73", X"6B", X"0D", X"0A", X"09", X"72", X"65", X"72", X"61", X"73", X"65", X"20", X"5B", X"70",
X"61", X"67", X"65", X"5D", X"09", X"09", X"09", X"45", X"72", X"61", X"73", X"65", X"20", X"52", X"41", X"4D",
X"20", X"64", X"69", X"73", X"6B", X"0D", X"0A", X"09", X"72", X"72", X"65", X"61", X"64", X"20", X"5B", X"70",
X"61", X"67", X"65", X"5D", X"20", X"5B", X"66", X"6C", X"61", X"73", X"68", X"70", X"61", X"67", X"65", X"5D",
X"09", X"52", X"65", X"61", X"64", X"20", X"52", X"41", X"4D", X"20", X"64", X"69", X"73", X"6B", X"20", X"66",
X"72", X"6F", X"6D", X"20", X"53", X"50", X"49", X"20", X"66", X"6C", X"61", X"73", X"68", X"0D", X"0A", X"09",
X"72", X"77", X"72", X"69", X"74", X"65", X"20", X"5B", X"70", X"61", X"67", X"65", X"5D", X"20", X"5B", X"66",
X"6C", X"61", X"73", X"68", X"70", X"61", X"67", X"65", X"5D", X"09", X"57", X"72", X"69", X"74", X"65", X"20",
X"52", X"41", X"4D", X"20", X"64", X"69", X"73", X"6B", X"20", X"74", X"6F", X"20", X"53", X"50", X"49", X"20",
X"66", X"6C", X"61", X"73", X"68", X"0D", X"0A", X"09", X"40", X"5B", X"63", X"6D", X"64", X"5D", X"09", X"09",
X"09", X"09", X"50", X"65", X"72", X"66", X"6F", X"72", X"6D", X"20", X"63", X"6F", X"6D", X"6D", X"61", X"6E",
X"64", X"20", X"77", X"69", X"74", X"68", X"6F", X"75", X"74", X"20", X"65", X"63", X"68", X"6F", X"20", X"6F",
X"72", X"20", X"74", X"65", X"72", X"6D", X"69", X"6E", X"61", X"6C", X"20", X"68", X"61", X"6E", X"64", X"6C",
X"69", X"6E", X"67", X"20", X"28", X"62", X"75", X"6C", X"6B", X"20", X"6F", X"70", X"65", X"72", X"61", X"74",
X"69", X"6F", X"6E", X"73", X"29", X"0D", X"0A", X"00", X"72", X"62", X"6F", X"6F", X"74", X"20", X"00", X"62",
X"75", X"66", X"00", X"63", X"70", X"20", X"00", X"64", X"6D", X"20", X"00", X"68", X"65", X"6C", X"70", X"00",
X"3F", X"00", X"69", X"6E", X"20", X"00", X"6D", X"6D", X"75", X"00", X"6F", X"75", X"74", X"20", X"00", X"72",
X"75", X"6E", X"20", X"00", X"73", X"70", X"00", X"77", X"6D", X"20", X"00", X"72", X"65", X"72", X"61", X"73",
X"65", X"00", X"72", X"72", X"65", X"61", X"64", X"00", X"72", X"77", X"72", X"69", X"74", X"65", X"00", X"23",
X"FD", X"D1", X"F2", X"27", X"FD", X"61", X"F1", X"2B", X"FD", X"E4", X"F0", X"30", X"FD", X"E4", X"F0", X"32",
X"FD", X"ED", X"F0", X"36", X"FD", X"18", X"F2", X"18", X"FD", X"B0", X"F1", X"3A", X"FD", X"15", X"F1", X"3F",
X"FD", X"A4", X"F1", X"47", X"FD", X"37", X"F1", X"44", X"FD", X"EE", X"F2", X"1F", X"FD", X"0F", X"F3", X"4B",
X"FD", X"2F", X"F3", X"52", X"FD", X"B5", X"F3", X"58", X"FD", X"6B", X"F4", X"00", X"00", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE",
X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE", X"FE"


     );

begin

  ram_process: process(clk, byte_rom)
  begin
      if rising_edge(clk) then
          -- latch the address, in order to infer a synchronous memory
          address_latch <= a;
      end if;
  end process;

  d <= byte_rom(to_integer(unsigned(address_latch)));

end arch;
